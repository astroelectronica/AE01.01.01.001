.title KiCad schematic
.include "models/C2012CH2W101J060AA_p.mod"
.include "models/C2012X7R2A104K125AA_p.mod"
.include "models/C2012X7R2E103K125AA_p.mod"
.include "models/ZXCT1080.spice.txt"
R1 /PWR_IN /PWR_OUT 0.1
R2 /PWR_IN /PWR_OUT 0.1
R3 /PWR_OUT /SN 10K
XU3 /PWR_IN /SN C2012CH2W101J060AA_p
XU2 +5V 0 C2012X7R2A104K125AA_p
R4 /OUT /VOCM 100
XU4 /OUT 0 C2012X7R2E103K125AA_p
XU1 0 +5V /PWR_IN /SN /VOCM ZXCT1080
V2 +5V 0 5
V1 /PWR_IN 0 {VIN}
I1 /PWR_OUT 0 {ILOAD}
.end
